library verilog;
use verilog.vl_types.all;
entity CompressionFunction_vlg_vec_tst is
end CompressionFunction_vlg_vec_tst;
